-- megafunction wizard: %RAM: 2-PORT%
-- GENERATION: STANDARD
-- VERSION: WM1.0
-- MODULE: altsyncram

-- ============================================================
-- File Name: g.vhd
-- Megafunction Name(s):
--          altsyncram
--
-- Simulation Library Files(s):
--          altera_mf
-- ============================================================
-- ************************************************************
-- THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
--
-- 11.1 Build 259 01/25/2012 SP 2 SJ Full Version
-- ************************************************************


--Copyright (C) 1991-2011 Altera Corporation
--Your use of Altera Corporation's design tools, logic functions
--and other software and tools, and its AMPP partner logic
--functions, and any output files from any of the foregoing
--(including device programming or simulation files), and any
--associated documentation or information are expressly subject
--to the terms and conditions of the Altera Program License
--Subscription Agreement, Altera MegaCore Function License
--Agreement, or other applicable license agreement, including,
--without limitation, that your use is for the sole purpose of
--programming logic devices manufactured by Altera and sold by
--Altera or its authorized distributors.  Please refer to the
--applicable agreement for further details.


--EDIT:

--DPRAM with the different Addresswith and Wordwith of Port A and B
--Byteenable at A
--No Register at the outputs

LIBRARY ieee;
USE ieee.std_logic_1164.all;

LIBRARY altera_mf;
USE altera_mf.all;

ENTITY DPRAM_Plus IS
    generic(gAddresswidthA:     natural :=7;
            gAddresswidthB:     natural :=6;
            gWordWidthA:        natural :=32;
            gWordWidthB:        natural :=64);
    PORT
    (
        address_a   : IN STD_LOGIC_VECTOR (gAddresswidthA-1 DOWNTO 0);
        address_b   : IN STD_LOGIC_VECTOR (gAddresswidthB-1 DOWNTO 0);
        byteena_a   : IN STD_LOGIC_VECTOR ((gWordWidthA/8)-1 DOWNTO 0) :=  (OTHERS => '1');
        byteena_b   : IN STD_LOGIC_VECTOR ((gWordWidthB/8)-1 DOWNTO 0) :=  (OTHERS => '1');
        clock_a     : IN STD_LOGIC  := '1';
        clock_b     : IN STD_LOGIC ;
        data_a      : IN STD_LOGIC_VECTOR (gWordWidthA-1 DOWNTO 0);
        data_b      : IN STD_LOGIC_VECTOR (gWordWidthB-1 DOWNTO 0);
        rden_a      : IN STD_LOGIC  := '1';
        rden_b      : IN STD_LOGIC  := '1';
        wren_a      : IN STD_LOGIC  := '0';
        wren_b      : IN STD_LOGIC  := '0';
        q_a         : OUT STD_LOGIC_VECTOR (gWordWidthA-1 DOWNTO 0);
        q_b         : OUT STD_LOGIC_VECTOR (gWordWidthB-1 DOWNTO 0)
    );
END DPRAM_Plus;


ARCHITECTURE SYN OF DPRAM_Plus IS

    SIGNAL sub_wire0    : STD_LOGIC_VECTOR (gWordWidthA-1 DOWNTO 0);
    SIGNAL sub_wire1    : STD_LOGIC_VECTOR (gWordWidthB-1 DOWNTO 0);



    COMPONENT altsyncram
    GENERIC (
        address_reg_b       : STRING;
        byte_size       : NATURAL;
        clock_enable_input_a        : STRING;
        clock_enable_input_b        : STRING;
        clock_enable_output_a       : STRING;
        clock_enable_output_b       : STRING;
        indata_reg_b        : STRING;
        intended_device_family      : STRING;
        lpm_type        : STRING;
        numwords_a      : NATURAL;
        numwords_b      : NATURAL;
        operation_mode      : STRING;
        outdata_aclr_a      : STRING;
        outdata_aclr_b      : STRING;
        outdata_reg_a       : STRING;
        outdata_reg_b       : STRING;
        power_up_uninitialized      : STRING;
        ram_block_type      : STRING;
        read_during_write_mode_port_a       : STRING;
        read_during_write_mode_port_b       : STRING;
        widthad_a       : NATURAL;
        widthad_b       : NATURAL;
        width_a     : NATURAL;
        width_b     : NATURAL;
        width_byteena_a     : NATURAL;
        width_byteena_b     : NATURAL;
        wrcontrol_wraddress_reg_b       : STRING
    );
    PORT (
            byteena_a   : IN STD_LOGIC_VECTOR ((gWordWidthA/8)-1 DOWNTO 0);
            byteena_b   : IN STD_LOGIC_VECTOR ((gWordWidthB/8)-1 DOWNTO 0);
            clock0  :   IN STD_LOGIC ;
            wren_a  :   IN STD_LOGIC ;
            rden_a  :   IN STD_LOGIC ;
            address_b:  IN STD_LOGIC_VECTOR (gAddresswidthB-1 DOWNTO 0);
            clock1  :   IN STD_LOGIC ;
            data_b  :   IN STD_LOGIC_VECTOR (gWordWidthB-1 DOWNTO 0);
            q_a :       OUT STD_LOGIC_VECTOR (gWordWidthA-1 DOWNTO 0);
            wren_b  :   IN STD_LOGIC ;
            rden_b  :   IN STD_LOGIC ;
            address_a:  IN STD_LOGIC_VECTOR (gAddresswidthA-1 DOWNTO 0);
            data_a  :   IN STD_LOGIC_VECTOR (gWordWidthA-1 DOWNTO 0);
            q_b :       OUT STD_LOGIC_VECTOR (gWordWidthB-1 DOWNTO 0)
    );
    END COMPONENT;

BEGIN
    q_a    <= sub_wire0(gWordWidthA-1 DOWNTO 0);
    q_b    <= sub_wire1(gWordWidthB-1 DOWNTO 0);

    altsyncram_component : altsyncram
    GENERIC MAP (
        address_reg_b => "CLOCK1",
        byte_size => 8,
        clock_enable_input_a => "BYPASS",
        clock_enable_input_b => "BYPASS",
        clock_enable_output_a => "BYPASS",
        clock_enable_output_b => "BYPASS",
        indata_reg_b => "CLOCK1",
        intended_device_family => "Cyclone IV E",
        lpm_type => "altsyncram",
        numwords_a => 2**gAddresswidthA,
        numwords_b => 2**gAddresswidthB,
        operation_mode => "BIDIR_DUAL_PORT",
        outdata_aclr_a => "NONE",
        outdata_aclr_b => "NONE",
        outdata_reg_a => "UNREGISTERED",
        outdata_reg_b => "UNREGISTERED",
        power_up_uninitialized => "FALSE",
        ram_block_type => "M9K",
        read_during_write_mode_port_a => "NEW_DATA_NO_NBE_READ",
        read_during_write_mode_port_b => "NEW_DATA_NO_NBE_READ",
        widthad_a => gAddresswidthA,
        widthad_b => gAddresswidthB,
        width_a => gWordWidthA,
        width_b => gWordWidthB,
        width_byteena_a => (gWordWidthA/8),
        width_byteena_b => (gWordWidthB/8),
        wrcontrol_wraddress_reg_b => "CLOCK1"
    )
    PORT MAP (
        byteena_a => byteena_a,
        byteena_b => byteena_b,
        clock0 => clock_a,
        wren_a => wren_a,
        clock1 => clock_b,
        rden_a => rden_a,
        wren_b => wren_b,
        address_a => address_a,
        data_a => data_a,
        rden_b => rden_b,
        address_b => address_b,
        data_b => data_b,
        q_a => sub_wire0,
        q_b => sub_wire1
    );



END SYN;

-- ============================================================
-- CNX file retrieval info
-- ============================================================
-- Retrieval info: PRIVATE: ADDRESSSTALL_A NUMERIC "0"
-- Retrieval info: PRIVATE: ADDRESSSTALL_B NUMERIC "0"
-- Retrieval info: PRIVATE: BYTEENA_ACLR_A NUMERIC "0"
-- Retrieval info: PRIVATE: BYTEENA_ACLR_B NUMERIC "0"
-- Retrieval info: PRIVATE: BYTE_ENABLE_A NUMERIC "0"
-- Retrieval info: PRIVATE: BYTE_ENABLE_B NUMERIC "0"
-- Retrieval info: PRIVATE: BYTE_SIZE NUMERIC "8"
-- Retrieval info: PRIVATE: BlankMemory NUMERIC "1"
-- Retrieval info: PRIVATE: CLOCK_ENABLE_INPUT_A NUMERIC "0"
-- Retrieval info: PRIVATE: CLOCK_ENABLE_INPUT_B NUMERIC "0"
-- Retrieval info: PRIVATE: CLOCK_ENABLE_OUTPUT_A NUMERIC "0"
-- Retrieval info: PRIVATE: CLOCK_ENABLE_OUTPUT_B NUMERIC "0"
-- Retrieval info: PRIVATE: CLRdata NUMERIC "0"
-- Retrieval info: PRIVATE: CLRq NUMERIC "0"
-- Retrieval info: PRIVATE: CLRrdaddress NUMERIC "0"
-- Retrieval info: PRIVATE: CLRrren NUMERIC "0"
-- Retrieval info: PRIVATE: CLRwraddress NUMERIC "0"
-- Retrieval info: PRIVATE: CLRwren NUMERIC "0"
-- Retrieval info: PRIVATE: Clock NUMERIC "5"
-- Retrieval info: PRIVATE: Clock_A NUMERIC "0"
-- Retrieval info: PRIVATE: Clock_B NUMERIC "0"
-- Retrieval info: PRIVATE: ECC NUMERIC "0"
-- Retrieval info: PRIVATE: ECC_PIPELINE_STAGE NUMERIC "0"
-- Retrieval info: PRIVATE: IMPLEMENT_IN_LES NUMERIC "0"
-- Retrieval info: PRIVATE: INDATA_ACLR_B NUMERIC "0"
-- Retrieval info: PRIVATE: INDATA_REG_B NUMERIC "1"
-- Retrieval info: PRIVATE: INIT_FILE_LAYOUT STRING "PORT_A"
-- Retrieval info: PRIVATE: INIT_TO_SIM_X NUMERIC "0"
-- Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Cyclone IV E"
-- Retrieval info: PRIVATE: JTAG_ENABLED NUMERIC "0"
-- Retrieval info: PRIVATE: JTAG_ID STRING "NONE"
-- Retrieval info: PRIVATE: MAXIMUM_DEPTH NUMERIC "0"
-- Retrieval info: PRIVATE: MEMSIZE NUMERIC "2048"
-- Retrieval info: PRIVATE: MEM_IN_BITS NUMERIC "0"
-- Retrieval info: PRIVATE: MIFfilename STRING ""
-- Retrieval info: PRIVATE: OPERATION_MODE NUMERIC "3"
-- Retrieval info: PRIVATE: OUTDATA_ACLR_B NUMERIC "0"
-- Retrieval info: PRIVATE: OUTDATA_REG_B NUMERIC "0"
-- Retrieval info: PRIVATE: RAM_BLOCK_TYPE NUMERIC "2"
-- Retrieval info: PRIVATE: READ_DURING_WRITE_MODE_MIXED_PORTS NUMERIC "2"
-- Retrieval info: PRIVATE: READ_DURING_WRITE_MODE_PORT_A NUMERIC "3"
-- Retrieval info: PRIVATE: READ_DURING_WRITE_MODE_PORT_B NUMERIC "3"
-- Retrieval info: PRIVATE: REGdata NUMERIC "1"
-- Retrieval info: PRIVATE: REGq NUMERIC "0"
-- Retrieval info: PRIVATE: REGrdaddress NUMERIC "0"
-- Retrieval info: PRIVATE: REGrren NUMERIC "0"
-- Retrieval info: PRIVATE: REGwraddress NUMERIC "1"
-- Retrieval info: PRIVATE: REGwren NUMERIC "1"
-- Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX STRING "0"
-- Retrieval info: PRIVATE: USE_DIFF_CLKEN NUMERIC "0"
-- Retrieval info: PRIVATE: UseDPRAM NUMERIC "1"
-- Retrieval info: PRIVATE: VarWidth NUMERIC "0"
-- Retrieval info: PRIVATE: WIDTH_READ_A NUMERIC "64"
-- Retrieval info: PRIVATE: WIDTH_READ_B NUMERIC "64"
-- Retrieval info: PRIVATE: WIDTH_WRITE_A NUMERIC "64"
-- Retrieval info: PRIVATE: WIDTH_WRITE_B NUMERIC "64"
-- Retrieval info: PRIVATE: WRADDR_ACLR_B NUMERIC "0"
-- Retrieval info: PRIVATE: WRADDR_REG_B NUMERIC "1"
-- Retrieval info: PRIVATE: WRCTRL_ACLR_B NUMERIC "0"
-- Retrieval info: PRIVATE: enable NUMERIC "0"
-- Retrieval info: PRIVATE: rden NUMERIC "0"
-- Retrieval info: LIBRARY: altera_mf altera_mf.altera_mf_components.all
-- Retrieval info: CONSTANT: ADDRESS_REG_B STRING "CLOCK1"
-- Retrieval info: CONSTANT: CLOCK_ENABLE_INPUT_A STRING "BYPASS"
-- Retrieval info: CONSTANT: CLOCK_ENABLE_INPUT_B STRING "BYPASS"
-- Retrieval info: CONSTANT: CLOCK_ENABLE_OUTPUT_A STRING "BYPASS"
-- Retrieval info: CONSTANT: CLOCK_ENABLE_OUTPUT_B STRING "BYPASS"
-- Retrieval info: CONSTANT: INDATA_REG_B STRING "CLOCK1"
-- Retrieval info: CONSTANT: INTENDED_DEVICE_FAMILY STRING "Cyclone IV E"
-- Retrieval info: CONSTANT: LPM_TYPE STRING "altsyncram"
-- Retrieval info: CONSTANT: NUMWORDS_A NUMERIC "32"
-- Retrieval info: CONSTANT: NUMWORDS_B NUMERIC "32"
-- Retrieval info: CONSTANT: OPERATION_MODE STRING "BIDIR_DUAL_PORT"
-- Retrieval info: CONSTANT: OUTDATA_ACLR_A STRING "NONE"
-- Retrieval info: CONSTANT: OUTDATA_ACLR_B STRING "NONE"
-- Retrieval info: CONSTANT: OUTDATA_REG_A STRING "UNREGISTERED"
-- Retrieval info: CONSTANT: OUTDATA_REG_B STRING "UNREGISTERED"
-- Retrieval info: CONSTANT: POWER_UP_UNINITIALIZED STRING "FALSE"
-- Retrieval info: CONSTANT: RAM_BLOCK_TYPE STRING "M9K"
-- Retrieval info: CONSTANT: READ_DURING_WRITE_MODE_PORT_A STRING "NEW_DATA_NO_NBE_READ"
-- Retrieval info: CONSTANT: READ_DURING_WRITE_MODE_PORT_B STRING "NEW_DATA_NO_NBE_READ"
-- Retrieval info: CONSTANT: WIDTHAD_A NUMERIC "5"
-- Retrieval info: CONSTANT: WIDTHAD_B NUMERIC "5"
-- Retrieval info: CONSTANT: WIDTH_A NUMERIC "64"
-- Retrieval info: CONSTANT: WIDTH_B NUMERIC "64"
-- Retrieval info: CONSTANT: WIDTH_BYTEENA_A NUMERIC "1"
-- Retrieval info: CONSTANT: WIDTH_BYTEENA_B NUMERIC "1"
-- Retrieval info: CONSTANT: WRCONTROL_WRADDRESS_REG_B STRING "CLOCK1"
-- Retrieval info: USED_PORT: address_a 0 0 5 0 INPUT NODEFVAL "address_a[4..0]"
-- Retrieval info: USED_PORT: address_b 0 0 5 0 INPUT NODEFVAL "address_b[4..0]"
-- Retrieval info: USED_PORT: clock_a 0 0 0 0 INPUT VCC "clock_a"
-- Retrieval info: USED_PORT: clock_b 0 0 0 0 INPUT NODEFVAL "clock_b"
-- Retrieval info: USED_PORT: data_a 0 0 64 0 INPUT NODEFVAL "data_a[63..0]"
-- Retrieval info: USED_PORT: data_b 0 0 64 0 INPUT NODEFVAL "data_b[63..0]"
-- Retrieval info: USED_PORT: q_a 0 0 64 0 OUTPUT NODEFVAL "q_a[63..0]"
-- Retrieval info: USED_PORT: q_b 0 0 64 0 OUTPUT NODEFVAL "q_b[63..0]"
-- Retrieval info: USED_PORT: wren_a 0 0 0 0 INPUT GND "wren_a"
-- Retrieval info: USED_PORT: wren_b 0 0 0 0 INPUT GND "wren_b"
-- Retrieval info: CONNECT: @address_a 0 0 5 0 address_a 0 0 5 0
-- Retrieval info: CONNECT: @address_b 0 0 5 0 address_b 0 0 5 0
-- Retrieval info: CONNECT: @clock0 0 0 0 0 clock_a 0 0 0 0
-- Retrieval info: CONNECT: @clock1 0 0 0 0 clock_b 0 0 0 0
-- Retrieval info: CONNECT: @data_a 0 0 64 0 data_a 0 0 64 0
-- Retrieval info: CONNECT: @data_b 0 0 64 0 data_b 0 0 64 0
-- Retrieval info: CONNECT: @wren_a 0 0 0 0 wren_a 0 0 0 0
-- Retrieval info: CONNECT: @wren_b 0 0 0 0 wren_b 0 0 0 0
-- Retrieval info: CONNECT: q_a 0 0 64 0 @q_a 0 0 64 0
-- Retrieval info: CONNECT: q_b 0 0 64 0 @q_b 0 0 64 0
-- Retrieval info: GEN_FILE: TYPE_NORMAL g.vhd TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL g.inc FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL g.cmp TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL g.bsf FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL g_inst.vhd FALSE
-- Retrieval info: LIB_FILE: altera_mf
